
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity nios_lights is
	port (
		clk        : in    std_logic;             
		leds     : out   std_logic_vector(3 downto 0); 
		reset  : in    std_logic;
		sdram_addr      : out   std_logic_vector(11 downto 0);  
		sdram_ba        : out   std_logic_vector(1 downto 0);  
		sdram_cas_n     : out   std_logic;                      
		sdram_cke       : out   std_logic;                    
		sdram_cs_n      : out   std_logic;                    
		sdram_dq        : inout std_logic_vector(31 downto 0);
		sdram_dqm       : out   std_logic_vector(3 downto 0); 
		sdram_ras_n     : out   std_logic;                                        
		sdram_we_n      : out   std_logic;                                        
		sdram_clk       : out   std_logic;                                        
		switches        : in    std_logic_vector(3 downto 0)
	);
end  nios_lights;

architecture rtl of nios_lights is
component lights is
	port (
		clk_clk         : in    std_logic                     := '0';             --       clk.clk
		leds_export     : out   std_logic_vector(3 downto 0);                     --      leds.export
		reset_reset_n   : in    std_logic                     := '0';             --     reset.reset_n
		sdram_addr      : out   std_logic_vector(11 downto 0);                    --     sdram.addr
		sdram_ba        : out   std_logic_vector(1 downto 0);                     --          .ba
		sdram_cas_n     : out   std_logic;                                        --          .cas_n
		sdram_cke       : out   std_logic;                                        --          .cke
		sdram_cs_n      : out   std_logic;                                        --          .cs_n
		sdram_dq        : inout std_logic_vector(31 downto 0) := (others => '0'); --          .dq
		sdram_dqm       : out   std_logic_vector(3 downto 0);                     --          .dqm
		sdram_ras_n     : out   std_logic;                                        --          .ras_n
		sdram_we_n      : out   std_logic;                                        --          .we_n
		sdram_clk_clk   : out   std_logic;                                        -- sdram_clk.clk
		switches_export : in    std_logic_vector(3 downto 0)  := (others => '0')  --  switches.export
	);
end component;

begin

NIOS:lights
port map(clk, leds,reset,sdram_addr,sdram_ba,sdram_cas_n,sdram_cke,sdram_cs_n,sdram_dq,sdram_dqm,sdram_ras_n,sdram_we_n,sdram_clk,switches);

end architecture rtl; -- of lights
