
module waves (
	clk_clk,
	reset_reset_n,
	sdram_clock_clk);	

	input		clk_clk;
	input		reset_reset_n;
	output		sdram_clock_clk;
endmodule
